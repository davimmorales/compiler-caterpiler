module simpleInstructionsRam(clock, address, iRAMOutput);
	 input [9:0] address;
	 input clock;
	 output [31:0] iRAMOutput;
	 integer firstClock = 0;
	 reg [31:0] instructionsRAM[240:0];

	 always @ ( posedge clock ) begin
	 	 if (firstClock==0) begin
 
	 	 instructionsRAM[0] = 32'b01011100000000000000000000000000;//Nop
	 	 instructionsRAM[1] = 32'b01001000000000000000000010010010;//Jump to #146
	 	 instructionsRAM[2] = 32'b01010000011000000000000000101010;//Load m[#42] to r[3]
	 	 instructionsRAM[3] = 32'b00000100011001110000000000000000;//ADDi r[3], #0 to r[7]
	 	 instructionsRAM[4] = 32'b01010100111000000000000000100111;//Store r[7] in m[#39]
	 	 instructionsRAM[5] = 32'b01010000011000000000000000101010;//Load m[#42] to r[3]
	 	 instructionsRAM[6] = 32'b00000100011001000000000000011011;//ADDi r[3], #27 to r[4]
	 	 instructionsRAM[7] = 32'b01110000100000010000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[8] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[9] = 32'b01010100111000000000000000101001;//Store r[7] in m[#41]
	 	 instructionsRAM[10] = 32'b01010000011000000000000000101010;//Load m[#42] to r[3]
	 	 instructionsRAM[11] = 32'b00000100011000010000000000000001;//ADDi r[3], #1 to r[1]
	 	 instructionsRAM[12] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[13] = 32'b01010100111000000000000000100110;//Store r[7] in m[#38]
	 	 instructionsRAM[14] = 32'b01010000011000000000000000100110;//Load m[#38] to r[3]
	 	 instructionsRAM[15] = 32'b01010000100000000000000000101000;//Load m[#40] to r[4]
	 	 instructionsRAM[16] = 32'b01001100011001000000100000000000;//SLT if r[3] < r[4], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[17] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[18] = 32'b00111100111000000000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[19] = 32'b01000000000000000000000000011000;//Branch on Zero #24
	 	 instructionsRAM[20] = 32'b01010000011000000000000000100110;//Load m[#38] to r[3]
	 	 instructionsRAM[21] = 32'b00000100011001000000000000011011;//ADDi r[3], #27 to r[4]
	 	 instructionsRAM[22] = 32'b01110000100000010000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[23] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[24] = 32'b00000100111000110000000000000000;//ADDi r[7], #0 to r[3]
	 	 instructionsRAM[25] = 32'b01010000100000000000000000101001;//Load m[#41] to r[4]
	 	 instructionsRAM[26] = 32'b01001100011001000000100000000000;//SLT if r[3] < r[4], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[27] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[28] = 32'b00111100111000000000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[29] = 32'b01000000000000000000000000001001;//Branch on Zero #9
	 	 instructionsRAM[30] = 32'b01010000011000000000000000100110;//Load m[#38] to r[3]
	 	 instructionsRAM[31] = 32'b00000100011001000000000000011011;//ADDi r[3], #27 to r[4]
	 	 instructionsRAM[32] = 32'b01110000100000010000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[33] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[34] = 32'b01010100111000000000000000101001;//Store r[7] in m[#41]
	 	 instructionsRAM[35] = 32'b01010000011000000000000000100110;//Load m[#38] to r[3]
	 	 instructionsRAM[36] = 32'b00000100011001110000000000000000;//ADDi r[3], #0 to r[7]
	 	 instructionsRAM[37] = 32'b01010100111000000000000000100111;//Store r[7] in m[#39]
	 	 instructionsRAM[38] = 32'b01010000011000000000000000100110;//Load m[#38] to r[3]
	 	 instructionsRAM[39] = 32'b00000100011000010000000000000001;//ADDi r[3], #1 to r[1]
	 	 instructionsRAM[40] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[41] = 32'b01010100111000000000000000100110;//Store r[7] in m[#38]
	 	 instructionsRAM[42] = 32'b01001000000000000000000000001110;//Jump to #14
	 	 instructionsRAM[43] = 32'b01010000001000000000000000100111;//Load m[#39] to r[1]
	 	 instructionsRAM[44] = 32'b00000100001111100000000000000000;//ADDi r[1], #0 to r[30]
	 	 instructionsRAM[45] = 32'b01110011111000010000000000000000;//Loadr m[r[31]] to r[1]
	 	 instructionsRAM[46] = 32'b01111000001000000000000000000000;//Jump to r[1]
	 	 instructionsRAM[47] = 32'b01110011111000010000000000000000;//Loadr m[r[31]] to r[1]
	 	 instructionsRAM[48] = 32'b01111000001000000000000000000000;//Jump to r[1]
	 	 instructionsRAM[49] = 32'b01010000011000000000000000011001;//Load m[#25] to r[3]
	 	 instructionsRAM[50] = 32'b00000100011001110000000000000000;//ADDi r[3], #0 to r[7]
	 	 instructionsRAM[51] = 32'b01010100111000000000000000010101;//Store r[7] in m[#21]
	 	 instructionsRAM[52] = 32'b01010000011000000000000000010111;//Load m[#23] to r[3]
	 	 instructionsRAM[53] = 32'b00001100011000010000000000000001;//SUBi r[3], #1 to r[1]
	 	 instructionsRAM[54] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[55] = 32'b01010000011000000000000000010101;//Load m[#21] to r[3]
	 	 instructionsRAM[56] = 32'b00000100111001000000000000000000;//ADDi r[7], #0 to r[4]
	 	 instructionsRAM[57] = 32'b01001100011001000000100000000000;//SLT if r[3] < r[4], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[58] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[59] = 32'b00111100111000000000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[60] = 32'b01000000000000000000000001010000;//Branch on Zero #80
	 	 instructionsRAM[61] = 32'b01010000001000000000000000001010;//Load m[#10] to r[1]
	 	 instructionsRAM[62] = 32'b01010000001000000000000000001010;//Load m[#10] to r[1]
	 	 instructionsRAM[63] = 32'b01010100001000000000000000011011;//Store r[1] in m[#27]
	 	 instructionsRAM[64] = 32'b01010000001000000000000000001011;//Load m[#11] to r[1]
	 	 instructionsRAM[65] = 32'b01010100001000000000000000011100;//Store r[1] in m[#28]
	 	 instructionsRAM[66] = 32'b01010000001000000000000000001100;//Load m[#12] to r[1]
	 	 instructionsRAM[67] = 32'b01010100001000000000000000011101;//Store r[1] in m[#29]
	 	 instructionsRAM[68] = 32'b01010000001000000000000000001101;//Load m[#13] to r[1]
	 	 instructionsRAM[69] = 32'b01010100001000000000000000011110;//Store r[1] in m[#30]
	 	 instructionsRAM[70] = 32'b01010000001000000000000000001110;//Load m[#14] to r[1]
	 	 instructionsRAM[71] = 32'b01010100001000000000000000011111;//Store r[1] in m[#31]
	 	 instructionsRAM[72] = 32'b01010000001000000000000000001111;//Load m[#15] to r[1]
	 	 instructionsRAM[73] = 32'b01010100001000000000000000100000;//Store r[1] in m[#32]
	 	 instructionsRAM[74] = 32'b01010000001000000000000000010000;//Load m[#16] to r[1]
	 	 instructionsRAM[75] = 32'b01010100001000000000000000100001;//Store r[1] in m[#33]
	 	 instructionsRAM[76] = 32'b01010000001000000000000000010001;//Load m[#17] to r[1]
	 	 instructionsRAM[77] = 32'b01010100001000000000000000100010;//Store r[1] in m[#34]
	 	 instructionsRAM[78] = 32'b01010000001000000000000000010010;//Load m[#18] to r[1]
	 	 instructionsRAM[79] = 32'b01010100001000000000000000100011;//Store r[1] in m[#35]
	 	 instructionsRAM[80] = 32'b01010000001000000000000000010011;//Load m[#19] to r[1]
	 	 instructionsRAM[81] = 32'b01010100001000000000000000100100;//Store r[1] in m[#36]
	 	 instructionsRAM[82] = 32'b01010000001000000000000000010100;//Load m[#20] to r[1]
	 	 instructionsRAM[83] = 32'b01010100001000000000000000100101;//Store r[1] in m[#37]
	 	 instructionsRAM[84] = 32'b01010000001000000000000000010101;//Load m[#21] to r[1]
	 	 instructionsRAM[85] = 32'b01010100001000000000000000101010;//Store r[1] in m[#42]
	 	 instructionsRAM[86] = 32'b01010000001000000000000000010111;//Load m[#23] to r[1]
	 	 instructionsRAM[87] = 32'b01010100001000000000000000101000;//Store r[1] in m[#40]
	 	 instructionsRAM[88] = 32'b01011011111000000000000000110111;//Loadi #55 to r[31]
	 	 instructionsRAM[89] = 32'b00000111111111110000000000000001;//ADDi r[31], #1 to r[31]
	 	 instructionsRAM[90] = 32'b01011000001000000000000001011101;//Loadi #93 to r[1]
	 	 instructionsRAM[91] = 32'b01110111111000010000000000000000;//Storer to r[1] in m[r[31]] 
	 	 instructionsRAM[92] = 32'b01001000000000000000000000000010;//Jump to #2
	 	 instructionsRAM[93] = 32'b00001111111111110000000000000001;//SUBi r[31], #1 to r[31]
	 	 instructionsRAM[94] = 32'b01010000001000000000000000011011;//Load m[#27] to r[1]
	 	 instructionsRAM[95] = 32'b01010100001000000000000000001010;//Store r[1] in m[#10]
	 	 instructionsRAM[96] = 32'b01010000001000000000000000011100;//Load m[#28] to r[1]
	 	 instructionsRAM[97] = 32'b01010100001000000000000000001011;//Store r[1] in m[#11]
	 	 instructionsRAM[98] = 32'b01010000001000000000000000011101;//Load m[#29] to r[1]
	 	 instructionsRAM[99] = 32'b01010100001000000000000000001100;//Store r[1] in m[#12]
	 	 instructionsRAM[100] = 32'b01010000001000000000000000011110;//Load m[#30] to r[1]
	 	 instructionsRAM[101] = 32'b01010100001000000000000000001101;//Store r[1] in m[#13]
	 	 instructionsRAM[102] = 32'b01010000001000000000000000011111;//Load m[#31] to r[1]
	 	 instructionsRAM[103] = 32'b01010100001000000000000000001110;//Store r[1] in m[#14]
	 	 instructionsRAM[104] = 32'b01010000001000000000000000100000;//Load m[#32] to r[1]
	 	 instructionsRAM[105] = 32'b01010100001000000000000000001111;//Store r[1] in m[#15]
	 	 instructionsRAM[106] = 32'b01010000001000000000000000100001;//Load m[#33] to r[1]
	 	 instructionsRAM[107] = 32'b01010100001000000000000000010000;//Store r[1] in m[#16]
	 	 instructionsRAM[108] = 32'b01010000001000000000000000100010;//Load m[#34] to r[1]
	 	 instructionsRAM[109] = 32'b01010100001000000000000000010001;//Store r[1] in m[#17]
	 	 instructionsRAM[110] = 32'b01010000001000000000000000100011;//Load m[#35] to r[1]
	 	 instructionsRAM[111] = 32'b01010100001000000000000000010010;//Store r[1] in m[#18]
	 	 instructionsRAM[112] = 32'b01010000001000000000000000100100;//Load m[#36] to r[1]
	 	 instructionsRAM[113] = 32'b01010100001000000000000000010011;//Store r[1] in m[#19]
	 	 instructionsRAM[114] = 32'b01010000001000000000000000100101;//Load m[#37] to r[1]
	 	 instructionsRAM[115] = 32'b01010100001000000000000000010100;//Store r[1] in m[#20]
	 	 instructionsRAM[116] = 32'b00000111110001110000000000000000;//ADDi r[30], #0 to r[7]
	 	 instructionsRAM[117] = 32'b01010100111000000000000000010110;//Store r[7] in m[#22]
	 	 instructionsRAM[118] = 32'b01010000011000000000000000010110;//Load m[#22] to r[3]
	 	 instructionsRAM[119] = 32'b00000100011001000000000000001010;//ADDi r[3], #10 to r[4]
	 	 instructionsRAM[120] = 32'b01110000100000010000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[121] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[122] = 32'b01010100111000000000000000011000;//Store r[7] in m[#24]
	 	 instructionsRAM[123] = 32'b01010000011000000000000000010101;//Load m[#21] to r[3]
	 	 instructionsRAM[124] = 32'b00000100011001000000000000001010;//ADDi r[3], #10 to r[4]
	 	 instructionsRAM[125] = 32'b01110000100000010000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[126] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[127] = 32'b01010000011000000000000000010110;//Load m[#22] to r[3]
	 	 instructionsRAM[128] = 32'b00000100011001000000000000001010;//ADDi r[3], #10 to r[4]
	 	 instructionsRAM[129] = 32'b01110100100001110000000000000000;//Storer to r[7] in m[r[4]] 
	 	 instructionsRAM[130] = 32'b01010000011000000000000000011000;//Load m[#24] to r[3]
	 	 instructionsRAM[131] = 32'b00000100011001110000000000000000;//ADDi r[3], #0 to r[7]
	 	 instructionsRAM[132] = 32'b01010000011000000000000000010101;//Load m[#21] to r[3]
	 	 instructionsRAM[133] = 32'b00000100011001000000000000001010;//ADDi r[3], #10 to r[4]
	 	 instructionsRAM[134] = 32'b01110100100001110000000000000000;//Storer to r[7] in m[r[4]] 
	 	 instructionsRAM[135] = 32'b01010000011000000000000000010101;//Load m[#21] to r[3]
	 	 instructionsRAM[136] = 32'b00000100011000010000000000000001;//ADDi r[3], #1 to r[1]
	 	 instructionsRAM[137] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[138] = 32'b01010100111000000000000000010101;//Store r[7] in m[#21]
	 	 instructionsRAM[139] = 32'b01001000000000000000000000110100;//Jump to #52
	 	 instructionsRAM[140] = 32'b01110011111000010000000000000000;//Loadr m[r[31]] to r[1]
	 	 instructionsRAM[141] = 32'b01111000001000000000000000000000;//Jump to r[1]
	 	 instructionsRAM[142] = 32'b01110011111000010000000000000000;//Loadr m[r[31]] to r[1]
	 	 instructionsRAM[143] = 32'b01111000001000000000000000000000;//Jump to r[1]
	 	 instructionsRAM[144] = 32'b01110011111000010000000000000000;//Loadr m[r[31]] to r[1]
	 	 instructionsRAM[145] = 32'b01111000001000000000000000000000;//Jump to r[1]
	 	 instructionsRAM[146] = 32'b01011000001000000000000000000000;//Loadi #0 to r[1]
	 	 instructionsRAM[147] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[148] = 32'b01010100111000000000000000001000;//Store r[7] in m[#8]
	 	 instructionsRAM[149] = 32'b01010000011000000000000000001000;//Load m[#8] to r[3]
	 	 instructionsRAM[150] = 32'b01011000100000000000000000001010;//Loadi #10 to r[4]
	 	 instructionsRAM[151] = 32'b01001100011001000000100000000000;//SLT if r[3] < r[4], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[152] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[153] = 32'b00111100111000000000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[154] = 32'b01000000000000000000000000001011;//Branch on Zero #11
	 	 instructionsRAM[155] = 32'b01100000001000000000000000000000;//Input to r[1]
	 	 instructionsRAM[156] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[157] = 32'b01010000011000000000000000001000;//Load m[#8] to r[3]
	 	 instructionsRAM[158] = 32'b00000100011001000000000000101100;//ADDi r[3], #44 to r[4]
	 	 instructionsRAM[159] = 32'b01110100100001110000000000000000;//Storer to r[7] in m[r[4]] 
	 	 instructionsRAM[160] = 32'b01010000011000000000000000001000;//Load m[#8] to r[3]
	 	 instructionsRAM[161] = 32'b00000100011000010000000000000001;//ADDi r[3], #1 to r[1]
	 	 instructionsRAM[162] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[163] = 32'b01010100111000000000000000001000;//Store r[7] in m[#8]
	 	 instructionsRAM[164] = 32'b01001000000000000000000010010101;//Jump to #149
	 	 instructionsRAM[165] = 32'b01010000001000000000000000101100;//Load m[#44] to r[1]
	 	 instructionsRAM[166] = 32'b01010000001000000000000000101100;//Load m[#44] to r[1]
	 	 instructionsRAM[167] = 32'b01010100001000000000000000001010;//Store r[1] in m[#10]
	 	 instructionsRAM[168] = 32'b01010000001000000000000000101101;//Load m[#45] to r[1]
	 	 instructionsRAM[169] = 32'b01010100001000000000000000001011;//Store r[1] in m[#11]
	 	 instructionsRAM[170] = 32'b01010000001000000000000000101110;//Load m[#46] to r[1]
	 	 instructionsRAM[171] = 32'b01010100001000000000000000001100;//Store r[1] in m[#12]
	 	 instructionsRAM[172] = 32'b01010000001000000000000000101111;//Load m[#47] to r[1]
	 	 instructionsRAM[173] = 32'b01010100001000000000000000001101;//Store r[1] in m[#13]
	 	 instructionsRAM[174] = 32'b01010000001000000000000000110000;//Load m[#48] to r[1]
	 	 instructionsRAM[175] = 32'b01010100001000000000000000001110;//Store r[1] in m[#14]
	 	 instructionsRAM[176] = 32'b01010000001000000000000000110001;//Load m[#49] to r[1]
	 	 instructionsRAM[177] = 32'b01010100001000000000000000001111;//Store r[1] in m[#15]
	 	 instructionsRAM[178] = 32'b01010000001000000000000000110010;//Load m[#50] to r[1]
	 	 instructionsRAM[179] = 32'b01010100001000000000000000010000;//Store r[1] in m[#16]
	 	 instructionsRAM[180] = 32'b01010000001000000000000000110011;//Load m[#51] to r[1]
	 	 instructionsRAM[181] = 32'b01010100001000000000000000010001;//Store r[1] in m[#17]
	 	 instructionsRAM[182] = 32'b01010000001000000000000000110100;//Load m[#52] to r[1]
	 	 instructionsRAM[183] = 32'b01010100001000000000000000010010;//Store r[1] in m[#18]
	 	 instructionsRAM[184] = 32'b01010000001000000000000000110101;//Load m[#53] to r[1]
	 	 instructionsRAM[185] = 32'b01010100001000000000000000010011;//Store r[1] in m[#19]
	 	 instructionsRAM[186] = 32'b01010000001000000000000000110110;//Load m[#54] to r[1]
	 	 instructionsRAM[187] = 32'b01010100001000000000000000010100;//Store r[1] in m[#20]
	 	 instructionsRAM[188] = 32'b01011000001000000000000000000000;//Loadi #0 to r[1]
	 	 instructionsRAM[189] = 32'b01010100001000000000000000011001;//Store r[1] in m[#25]
	 	 instructionsRAM[190] = 32'b01011000001000000000000000001010;//Loadi #10 to r[1]
	 	 instructionsRAM[191] = 32'b01010100001000000000000000010111;//Store r[1] in m[#23]
	 	 instructionsRAM[192] = 32'b00000111111111110000000000000001;//ADDi r[31], #1 to r[31]
	 	 instructionsRAM[193] = 32'b01011000001000000000000011000100;//Loadi #196 to r[1]
	 	 instructionsRAM[194] = 32'b01110111111000010000000000000000;//Storer to r[1] in m[r[31]] 
	 	 instructionsRAM[195] = 32'b01001000000000000000000000110001;//Jump to #49
	 	 instructionsRAM[196] = 32'b00001111111111110000000000000001;//SUBi r[31], #1 to r[31]
	 	 instructionsRAM[197] = 32'b01010000001000000000000000001010;//Load m[#10] to r[1]
	 	 instructionsRAM[198] = 32'b01010100001000000000000000101100;//Store r[1] in m[#44]
	 	 instructionsRAM[199] = 32'b01010000001000000000000000001011;//Load m[#11] to r[1]
	 	 instructionsRAM[200] = 32'b01010100001000000000000000101101;//Store r[1] in m[#45]
	 	 instructionsRAM[201] = 32'b01010000001000000000000000001100;//Load m[#12] to r[1]
	 	 instructionsRAM[202] = 32'b01010100001000000000000000101110;//Store r[1] in m[#46]
	 	 instructionsRAM[203] = 32'b01010000001000000000000000001101;//Load m[#13] to r[1]
	 	 instructionsRAM[204] = 32'b01010100001000000000000000101111;//Store r[1] in m[#47]
	 	 instructionsRAM[205] = 32'b01010000001000000000000000001110;//Load m[#14] to r[1]
	 	 instructionsRAM[206] = 32'b01010100001000000000000000110000;//Store r[1] in m[#48]
	 	 instructionsRAM[207] = 32'b01010000001000000000000000001111;//Load m[#15] to r[1]
	 	 instructionsRAM[208] = 32'b01010100001000000000000000110001;//Store r[1] in m[#49]
	 	 instructionsRAM[209] = 32'b01010000001000000000000000010000;//Load m[#16] to r[1]
	 	 instructionsRAM[210] = 32'b01010100001000000000000000110010;//Store r[1] in m[#50]
	 	 instructionsRAM[211] = 32'b01010000001000000000000000010001;//Load m[#17] to r[1]
	 	 instructionsRAM[212] = 32'b01010100001000000000000000110011;//Store r[1] in m[#51]
	 	 instructionsRAM[213] = 32'b01010000001000000000000000010010;//Load m[#18] to r[1]
	 	 instructionsRAM[214] = 32'b01010100001000000000000000110100;//Store r[1] in m[#52]
	 	 instructionsRAM[215] = 32'b01010000001000000000000000010011;//Load m[#19] to r[1]
	 	 instructionsRAM[216] = 32'b01010100001000000000000000110101;//Store r[1] in m[#53]
	 	 instructionsRAM[217] = 32'b01010000001000000000000000010100;//Load m[#20] to r[1]
	 	 instructionsRAM[218] = 32'b01010100001000000000000000110110;//Store r[1] in m[#54]
	 	 instructionsRAM[219] = 32'b01011000001000000000000000000000;//Loadi #0 to r[1]
	 	 instructionsRAM[220] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[221] = 32'b01010100111000000000000000001000;//Store r[7] in m[#8]
	 	 instructionsRAM[222] = 32'b01010000011000000000000000001000;//Load m[#8] to r[3]
	 	 instructionsRAM[223] = 32'b01011000100000000000000000001010;//Loadi #10 to r[4]
	 	 instructionsRAM[224] = 32'b01001100011001000000100000000000;//SLT if r[3] < r[4], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[225] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[226] = 32'b00111100111000000000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[227] = 32'b01000000000000000000000000001101;//Branch on Zero #13
	 	 instructionsRAM[228] = 32'b01010000011000000000000000001000;//Load m[#8] to r[3]
	 	 instructionsRAM[229] = 32'b00000100011001000000000000101100;//ADDi r[3], #44 to r[4]
	 	 instructionsRAM[230] = 32'b01110000100000010000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[231] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[232] = 32'b00000100111000010000000000000000;//ADDi r[7], #0 to r[1]
	 	 instructionsRAM[233] = 32'b01101000001000000000000000000000;//Pre Output r[1]
	 	 instructionsRAM[234] = 32'b01101100001000000000000000000000;//Output r[1]
	 	 instructionsRAM[235] = 32'b01010000011000000000000000001000;//Load m[#8] to r[3]
	 	 instructionsRAM[236] = 32'b00000100011000010000000000000001;//ADDi r[3], #1 to r[1]
	 	 instructionsRAM[237] = 32'b00000100001001110000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[238] = 32'b01010100111000000000000000001000;//Store r[7] in m[#8]
	 	 instructionsRAM[239] = 32'b01001000000000000000000011011110;//Jump to #222

	 	 firstClock <= 0;
	 	 end
	 end

	 assign iRAMOutput = instructionsRAM[address];
endmodule // simpleInstructionsRAM
