module simpleInstructionsRam(clock, address, iRAMOutput);
	 input [9:0] address;
	 input clock;
	 output [31:0] iRAMOutput;
	 integer firstClock = 0;
	 reg [31:0] instructionsRAM[159:0];

	 always @ ( posedge clock ) begin
	 	 if (firstClock==0) begin
 
	 	 instructionsRAM[0] = 32'b01101100000000000000000000000000;//Nop
	 	 instructionsRAM[1] = 32'b01010100000000000000000001010100;//Jump to #84
	 	 instructionsRAM[2] = 32'b01101000001000000000000000000100;//Loadi #4 to r[1]
	 	 instructionsRAM[3] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[4] = 32'b01100100111000000000000000000010;//Store r[7] in m[#2]
	 	 instructionsRAM[5] = 32'b01100000001000000000000000000010;//Load m[#2] to r[1]
	 	 instructionsRAM[6] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[7] = 32'b01100000011000000000000000000010;//Load m[#2] to r[3]
	 	 instructionsRAM[8] = 32'b01101000100000000000000000000000;//Loadi #0 to r[4]
	 	 instructionsRAM[9] = 32'b01011100001001000001100000000000;//SLT if r[4] < r[3], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[10] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[11] = 32'b01111100000001110000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[12] = 32'b01001100000000000000000001000101;//Branch on Zero #69
	 	 instructionsRAM[13] = 32'b01101000001000000000000000000000;//Loadi #0 to r[1]
	 	 instructionsRAM[14] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[15] = 32'b01100100111000000000000000000001;//Store r[7] in m[#1]
	 	 instructionsRAM[16] = 32'b01100000011000000000000000000001;//Load m[#1] to r[3]
	 	 instructionsRAM[17] = 32'b01100000100000000000000000000010;//Load m[#2] to r[4]
	 	 instructionsRAM[18] = 32'b01011100001000110010000000000000;//SLT if r[3] < r[4], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[19] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[20] = 32'b01111100000001110000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[21] = 32'b01001100000000000000000000110111;//Branch on Zero #55
	 	 instructionsRAM[22] = 32'b01100000011000000000000000000001;//Load m[#1] to r[3]
	 	 instructionsRAM[23] = 32'b00000100001000110000000000000001;//ADDi r[3], #1 to r[1]
	 	 instructionsRAM[24] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[25] = 32'b01100100111000000000000000000011;//Store r[7] in m[#3]
	 	 instructionsRAM[26] = 32'b01100000011000000000000000000001;//Load m[#1] to r[3]
	 	 instructionsRAM[27] = 32'b00000100100000110000000000000101;//ADDi r[3], #5 to r[4]
	 	 instructionsRAM[28] = 32'b10000100001001000000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[29] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[30] = 32'b01100000011000000000000000000011;//Load m[#3] to r[3]
	 	 instructionsRAM[31] = 32'b00000100100000110000000000000101;//ADDi r[3], #5 to r[4]
	 	 instructionsRAM[32] = 32'b10000100001001000000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[33] = 32'b00000101000000010000000000000000;//ADDi r[1], #0 to r[8]
	 	 instructionsRAM[34] = 32'b00000100011001110000000000000000;//ADDi r[7], #0 to r[3]
	 	 instructionsRAM[35] = 32'b00000100100010000000000000000000;//ADDi r[8], #0 to r[4]
	 	 instructionsRAM[36] = 32'b01011100001001000001100000000000;//SLT if r[4] < r[3], r[1] = 1 else r[1] = 0
	 	 instructionsRAM[37] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[38] = 32'b01111100000001110000000000000000;//Pre Branch r[7]
	 	 instructionsRAM[39] = 32'b01001100000000000000000000100000;//Branch on Zero #32
	 	 instructionsRAM[40] = 32'b01100000001000000000000000000001;//Load m[#1] to r[1]
	 	 instructionsRAM[41] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[42] = 32'b01100000001000000000000000000011;//Load m[#3] to r[1]
	 	 instructionsRAM[43] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[44] = 32'b01100000001000000000000000000010;//Load m[#2] to r[1]
	 	 instructionsRAM[45] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[46] = 32'b01100000011000000000000000000001;//Load m[#1] to r[3]
	 	 instructionsRAM[47] = 32'b00000100100000110000000000000101;//ADDi r[3], #5 to r[4]
	 	 instructionsRAM[48] = 32'b10000100001001000000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[49] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[50] = 32'b01100100111000000000000000001011;//Store r[7] in m[#11]
	 	 instructionsRAM[51] = 32'b01100000011000000000000000000011;//Load m[#3] to r[3]
	 	 instructionsRAM[52] = 32'b00000100100000110000000000000101;//ADDi r[3], #5 to r[4]
	 	 instructionsRAM[53] = 32'b10000100001001000000000000000000;//Loadr m[r[4]] to r[1]
	 	 instructionsRAM[54] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[55] = 32'b01100100111000000000000000001100;//Store r[7] in m[#12]
	 	 instructionsRAM[56] = 32'b01100000011000000000000000001100;//Load m[#12] to r[3]
	 	 instructionsRAM[57] = 32'b00000100111000110000000000000000;//ADDi r[3], #0 to r[7]
	 	 instructionsRAM[58] = 32'b01100000011000000000000000000001;//Load m[#1] to r[3]
	 	 instructionsRAM[59] = 32'b00000100100000110000000000000101;//ADDi r[3], #5 to r[4]
	 	 instructionsRAM[60] = 32'b10001000111001000000000000000000;//rStore to r[7] in m[r[4]] 
	 	 instructionsRAM[61] = 32'b01100000011000000000000000001011;//Load m[#11] to r[3]
	 	 instructionsRAM[62] = 32'b00000100111000110000000000000000;//ADDi r[3], #0 to r[7]
	 	 instructionsRAM[63] = 32'b01100000011000000000000000000011;//Load m[#3] to r[3]
	 	 instructionsRAM[64] = 32'b00000100100000110000000000000101;//ADDi r[3], #5 to r[4]
	 	 instructionsRAM[65] = 32'b10001000111001000000000000000000;//rStore to r[7] in m[r[4]] 
	 	 instructionsRAM[66] = 32'b01100000001000000000000000000001;//Load m[#1] to r[1]
	 	 instructionsRAM[67] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[68] = 32'b01100000001000000000000000000011;//Load m[#3] to r[1]
	 	 instructionsRAM[69] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[70] = 32'b01100000001000000000000000000010;//Load m[#2] to r[1]
	 	 instructionsRAM[71] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[72] = 32'b01100000011000000000000000000001;//Load m[#1] to r[3]
	 	 instructionsRAM[73] = 32'b00000100001000110000000000000001;//ADDi r[3], #1 to r[1]
	 	 instructionsRAM[74] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[75] = 32'b01100100111000000000000000000001;//Store r[7] in m[#1]
	 	 instructionsRAM[76] = 32'b01010100000000000000000000010000;//Jump to #16
	 	 instructionsRAM[77] = 32'b01100000011000000000000000000010;//Load m[#2] to r[3]
	 	 instructionsRAM[78] = 32'b00001100001000110000000000000001;//SUBi r[3], #1 to r[1]
	 	 instructionsRAM[79] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[80] = 32'b01100100111000000000000000000010;//Store r[7] in m[#2]
	 	 instructionsRAM[81] = 32'b01010100000000000000000000000111;//Jump to #7
	 	 instructionsRAM[82] = 32'b10000100001111110000000000000000;//Loadr m[r[31]] to r[1]
	 	 instructionsRAM[83] = 32'b10001100000000010000000000000000;//Jump to r[1]
	 	 instructionsRAM[84] = 32'b01101000001000000000000000001111;//Loadi #15 to r[1]
	 	 instructionsRAM[85] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[86] = 32'b01100100111000000000000000010000;//Store r[7] in m[#16]
	 	 instructionsRAM[87] = 32'b01101000001000000000000001001000;//Loadi #72 to r[1]
	 	 instructionsRAM[88] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[89] = 32'b01100100111000000000000000010001;//Store r[7] in m[#17]
	 	 instructionsRAM[90] = 32'b01101000001000000000000000001110;//Loadi #14 to r[1]
	 	 instructionsRAM[91] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[92] = 32'b01100100111000000000000000010010;//Store r[7] in m[#18]
	 	 instructionsRAM[93] = 32'b01101000001000000000000000000001;//Loadi #1 to r[1]
	 	 instructionsRAM[94] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[95] = 32'b01100100111000000000000000010011;//Store r[7] in m[#19]
	 	 instructionsRAM[96] = 32'b01101000001000000000000000000011;//Loadi #3 to r[1]
	 	 instructionsRAM[97] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[98] = 32'b01100100111000000000000000010100;//Store r[7] in m[#20]
	 	 instructionsRAM[99] = 32'b01101000001000000000000000000101;//Loadi #5 to r[1]
	 	 instructionsRAM[100] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[101] = 32'b01100100111000000000000000010110;//Store r[7] in m[#22]
	 	 instructionsRAM[102] = 32'b01100000001000000000000000010000;//Load m[#16] to r[1]
	 	 instructionsRAM[103] = 32'b01100000001000000000000000010000;//Load m[#16] to r[1]
	 	 instructionsRAM[104] = 32'b01100100001000000000000000000101;//Store r[1] in m[#5]
	 	 instructionsRAM[105] = 32'b01100000001000000000000000010001;//Load m[#17] to r[1]
	 	 instructionsRAM[106] = 32'b01100100001000000000000000000110;//Store r[1] in m[#6]
	 	 instructionsRAM[107] = 32'b01100000001000000000000000010010;//Load m[#18] to r[1]
	 	 instructionsRAM[108] = 32'b01100100001000000000000000000111;//Store r[1] in m[#7]
	 	 instructionsRAM[109] = 32'b01100000001000000000000000010011;//Load m[#19] to r[1]
	 	 instructionsRAM[110] = 32'b01100100001000000000000000001000;//Store r[1] in m[#8]
	 	 instructionsRAM[111] = 32'b01100000001000000000000000010100;//Load m[#20] to r[1]
	 	 instructionsRAM[112] = 32'b01100100001000000000000000001001;//Store r[1] in m[#9]
	 	 instructionsRAM[113] = 32'b01100000001000000000000000010101;//Load m[#21] to r[1]
	 	 instructionsRAM[114] = 32'b01100100001000000000000000001010;//Store r[1] in m[#10]
	 	 instructionsRAM[115] = 32'b01100000001000000000000000010110;//Load m[#22] to r[1]
	 	 instructionsRAM[116] = 32'b01100100001000000000000000000000;//Store r[1] in m[#0]
	 	 instructionsRAM[117] = 32'b01101011111000000000000000011001;//Loadi #25 to r[31]
	 	 instructionsRAM[118] = 32'b00000111111111110000000000000001;//ADDi r[31], #1 to r[31]
	 	 instructionsRAM[119] = 32'b01101000001000000000000001111010;//Loadi #122 to r[1]
	 	 instructionsRAM[120] = 32'b10001000001111110000000000000000;//rStore to r[1] in m[r[31]] 
	 	 instructionsRAM[121] = 32'b01010100000000000000000000000010;//Jump to #2
	 	 instructionsRAM[122] = 32'b00001111111111110000000000000001;//SUBi r[31], #1 to r[31]
	 	 instructionsRAM[123] = 32'b01100000001000000000000000000101;//Load m[#5] to r[1]
	 	 instructionsRAM[124] = 32'b01100100001000000000000000010000;//Store r[1] in m[#16]
	 	 instructionsRAM[125] = 32'b01100000001000000000000000000110;//Load m[#6] to r[1]
	 	 instructionsRAM[126] = 32'b01100100001000000000000000010001;//Store r[1] in m[#17]
	 	 instructionsRAM[127] = 32'b01100000001000000000000000000111;//Load m[#7] to r[1]
	 	 instructionsRAM[128] = 32'b01100100001000000000000000010010;//Store r[1] in m[#18]
	 	 instructionsRAM[129] = 32'b01100000001000000000000000001000;//Load m[#8] to r[1]
	 	 instructionsRAM[130] = 32'b01100100001000000000000000010011;//Store r[1] in m[#19]
	 	 instructionsRAM[131] = 32'b01100000001000000000000000001001;//Load m[#9] to r[1]
	 	 instructionsRAM[132] = 32'b01100100001000000000000000010100;//Store r[1] in m[#20]
	 	 instructionsRAM[133] = 32'b01100000001000000000000000001010;//Load m[#10] to r[1]
	 	 instructionsRAM[134] = 32'b01100100001000000000000000010101;//Store r[1] in m[#21]
	 	 instructionsRAM[135] = 32'b01101000001000000000000000000000;//Loadi #0 to r[1]
	 	 instructionsRAM[136] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[137] = 32'b01100100111000000000000000010111;//Store r[7] in m[#23]
	 	 instructionsRAM[138] = 32'b01100000001000000000000000010000;//Load m[#16] to r[1]
	 	 instructionsRAM[139] = 32'b00000100111000010000000000000000;//ADDi r[1], #0 to r[7]
	 	 instructionsRAM[140] = 32'b00000100001001110000000000000000;//ADDi r[7], #0 to r[1]
	 	 instructionsRAM[141] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[142] = 32'b01100000001000000000000000010001;//Load m[#17] to r[1]
	 	 instructionsRAM[143] = 32'b00000101000000010000000000000000;//ADDi r[1], #0 to r[8]
	 	 instructionsRAM[144] = 32'b00000100001010000000000000000000;//ADDi r[8], #0 to r[1]
	 	 instructionsRAM[145] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[146] = 32'b01100000001000000000000000010010;//Load m[#18] to r[1]
	 	 instructionsRAM[147] = 32'b00000101001000010000000000000000;//ADDi r[1], #0 to r[9]
	 	 instructionsRAM[148] = 32'b00000100001010010000000000000000;//ADDi r[9], #0 to r[1]
	 	 instructionsRAM[149] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[150] = 32'b01100000001000000000000000010011;//Load m[#19] to r[1]
	 	 instructionsRAM[151] = 32'b00000101010000010000000000000000;//ADDi r[1], #0 to r[10]
	 	 instructionsRAM[152] = 32'b00000100001010100000000000000000;//ADDi r[10], #0 to r[1]
	 	 instructionsRAM[153] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[154] = 32'b01100000001000000000000000010100;//Load m[#20] to r[1]
	 	 instructionsRAM[155] = 32'b00000101011000010000000000000000;//ADDi r[1], #0 to r[11]
	 	 instructionsRAM[156] = 32'b00000100001010110000000000000000;//ADDi r[11], #0 to r[1]
	 	 instructionsRAM[157] = 32'b10000000001000000000000000000000;//Output r[1]
	 	 instructionsRAM[158] = 32'b01110000000000000000000000000000;//Hlt

	 	 firstClock <= 0;
	 	 end
	 end

	 assign iRAMOutput = instructionsRAM[address];
endmodule // simpleInstructionsRAM
